/*
	CEFET-MG
	Disciplina de Laboratório de Arquitetura e Organização de Computadores
	Data: 28/08/2021
	Aluno: Fernando Veizaga
	Matricula: 20203001902
*/

module extensor1p3(entrada, saida);
	input entrada;
	
	output reg [2:0] saida;
	
	always @ (entrada)
	begin
		saida <= {{2{1'b0}}, entrada};
	end
endmodule


module test_extensor1p3;
	reg ent;
	
	wire [2:0] saida;
	
	initial begin
		ent = 0;
		#2 ent = 1;
		#2 ent = 0;
	end
	
	initial begin
 		$monitor("Time=%0d entrada=%b saida=%b",$time, ent, saida);
 	end
	
	extensor1p3 mod1(ent, saida);
	
endmodule
